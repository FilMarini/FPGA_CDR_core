../locker_manager.vhd