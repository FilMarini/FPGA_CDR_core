../phase_detector.vhd