../phase_detector_unit/phase_detector.vhd