../top_level.vhd