../BBPFD.vhd