../slow_clock_pulse.vhd