../n_cycle_stuff/n_cycle_generator.vhd