../locker_monitoring.vhd