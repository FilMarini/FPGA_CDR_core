../PRBSpack.vhd