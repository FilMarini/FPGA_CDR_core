../frequency_detector_unit/quadrant_detector.vhd