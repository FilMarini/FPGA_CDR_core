../n_cycle_generator.vhd