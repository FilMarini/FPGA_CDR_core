../../GCU_utils.vhd