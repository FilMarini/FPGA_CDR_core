../phase_detector_unit/freq_controller.vhd