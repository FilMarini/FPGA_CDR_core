../n_cycle_stuff/n_cycle_calc.vhd