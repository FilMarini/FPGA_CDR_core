../n_cycle_stuff/slow_phase_analyzer.vhd