../GCU_utils.vhd