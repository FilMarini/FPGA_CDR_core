../n_cycle_stuff/deglitcher.vhd