../prbs_any.vhd