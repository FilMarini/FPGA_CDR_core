../clk_wiz.vhd