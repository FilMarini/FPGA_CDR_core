-------------------------------------------------------------------------------
-- Title      : Testbench for design "BBPD"
-- Project    : 
-------------------------------------------------------------------------------
-- File       : BBPD_tb.vhd
-- Author     : Filippo Marini   <filippo.marini@pd.infn.it>
-- Company    : Universita degli studi di Padova
-- Created    : 2019-12-09
-- Last update: 2019-12-09
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2019 Universita degli studi di Padova
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2019-12-09  1.0      filippo	Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

-------------------------------------------------------------------------------

entity BBPD_tb is

end entity BBPD_tb;

-------------------------------------------------------------------------------

architecture beh of BBPD_tb is

  -- component ports
  signal data_i    : std_logic;
  signal pd_o      : std_logic;

  -- clock
  signal clk_i : std_logic := '1';
  signal clk_180_i : std_logic := '0';

begin  -- architecture beh

  -- component instantiation
  DUT: entity work.BBPD
    port map (
      clk_i     => clk_i,
      clk_180_i => clk_180_i,
      data_i    => data_i,
      pd_o      => pd_o);

  -- clock generation
  clk_i <= not clk_i after 8 ns;
  clk_180_i <= not clk_180_i after 8 ns;

  -- waveform generation
  WaveGen_Proc: process
  begin
    data_i <= '0';
    wait for 1 ns;  -- insert signal assignments here
    while true loop
      data_i <= '0';
      wait for 16 ns;
      data_i <= '1';
      wait for 16 ns;
      data_i <= '0';
      wait for 16 ns;
      data_i <= '1';
      wait for 16 ns;
      data_i <= '1';
      wait for 16 ns;
      data_i <= '0';
      wait for 16 ns;
      data_i <= '1';
      wait for 16 ns;
      data_i <= '0';
      wait for 16 ns;
      data_i <= '1';
      wait for 16 ns;
      data_i <= '0';
      wait for 16 ns;
      data_i <= '1';
    end loop;
    wait;
    
  end process WaveGen_Proc;

  

end architecture beh;

-------------------------------------------------------------------------------

-- configuration BBPD_tb_beh_cfg of BBPD_tb is
--   for beh
--   end for;
-- end BBPD_tb_beh_cfg;

-------------------------------------------------------------------------------
