../frequency_detector.vhd