../pfd.vhd