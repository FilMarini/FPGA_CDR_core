../deglitcher.vhd