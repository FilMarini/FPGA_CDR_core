../phase_detector_unit/phase_shift_filter_slave.vhd