../lock_manager.vhd