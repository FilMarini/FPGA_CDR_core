../BBPD.vhd