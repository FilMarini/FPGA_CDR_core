../frequency_detector_unit/quadrant_shifting_detector.vhd